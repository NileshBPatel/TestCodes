program hello;
  
  inital begin
    $display("HelloWorld");    
  end

endprogram 
